`define DSP_PORT_SIZE_A 24
`define DSP_PORT_SIZE_B 17