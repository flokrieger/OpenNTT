/*
    OpenNTT - 2024
    Florian Krieger, Florian Hirner, Ahmet Can Mert, Sujoy Sinha Roy
    Contact: florian.krieger@iaik.tugraz.at
*/

package intmul_pkg;
  localparam DSP_PORT_SIZE_A = 24;
  localparam DSP_PORT_SIZE_B = 17;
endpackage